`timescale 1ns / 1ps
`include "mycpu.svh"
module hazard(
    //from ID_STAGE

    //to ID_STAGE


    //from EXE_STAGE


    //from  MEM_STAGE 单元


    //from WB_STAGE

);

//**********************//********************//
    //阻塞逻辑设计
    // 1. LW阻塞检测

    // 2. 分支阻塞检测

    // 3. 阻塞结果输出

//**********************//********************//

//**********************//********************//
    // 前递设计包括
    // 1 LW引起的阻塞检测

    //2 前递逻辑判断

    //3 前递结果输出

//********************//******************//
 
endmodule
