/*------------------------------------------------------------------------------
--------------------------------------------------------------------------------
Copyright (c) 2016, Loongson Technology Corporation Limited.

All rights reserved.

Redistribution and use in source and binary forms, with or without modification,
are permitted provided that the following conditions are met:

1. Redistributions of source code must retain the above copyright notice, this 
list of conditions and the following disclaimer.

2. Redistributions in binary form must reproduce the above copyright notice, 
this list of conditions and the following disclaimer in the documentation and/or
other materials provided with the distribution.

3. Neither the name of Loongson Technology Corporation Limited nor the names of 
its contributors may be used to endorse or promote products derived from this 
software without specific prior written permission.

THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND 
ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED 
WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE 
DISCLAIMED. IN NO EVENT SHALL LOONGSON TECHNOLOGY CORPORATION LIMITED BE LIABLE
TO ANY PARTY FOR DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR 
CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE 
GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) 
HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT 
LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF
THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
--------------------------------------------------------------------------------
------------------------------------------------------------------------------*/

//*************************************************************************
//   > File Name   : soc_mini_top.v
//   > Description : SoC, included cpu, 
//                   inst ram, confreg
// 
//           -------------------------
//           |           cpu         |
//           -------------------------
//         inst|                  | data
//             |                  | 
//             |                  |           
//             |                  |           
//      -------------         -----------
//      | inst ram  |         | confreg |
//      -------------         -----------
//
//   > Author      : LOONGSON
//   > Date        : 2017-08-04
//*************************************************************************
`timescale 1ns / 1ps
`include "async_ram.sv"
`include "../mycpu/minicpu_top.sv"
`default_nettype none

//for simulation:
//1. if define SIMU_USE_PLL = 1, will use clk_pll to generate cpu_clk,
//   and simulation will be very slow.
//2. usually, please define SIMU_USE_PLL=0 to speed up simulation by assign
//   cpu_clk = clk.
//   at this time, cpu_clk frequency are both 100MHz, same as clk.
`define SIMU_USE_PLL 0 //set 0 to speed up simulation

module soc_mini_top #(parameter SIMULATION=1'b0)
(
    input          resetn, 
    input          clk,

    //------gpio-------
    output  [15:0] led,
    input   [7 :0] switch_1 
);

//clk and resetn
logic cpu_clk;
logic cpu_resetn;
always @(posedge cpu_clk)
begin
    cpu_resetn <= resetn;
end
assign cpu_clk   = clk;
// generate if(SIMULATION && `SIMU_USE_PLL==0)
// begin: speedup_simulation
//     assign cpu_clk   = clk;
// end
// else
// begin: pll
//     clk_pll clk_pll
//     (
//         .clk_in1 (clk),
//         .cpu_clk (cpu_clk),
//         .timer_clk ()
//     );
// end
// endgenerate

//cpu inst sram
logic        cpu_inst_we;
logic [31:0] cpu_inst_addr;
logic [31:0] cpu_inst_wdata;
logic [31:0] cpu_inst_rdata;
//cpu data sram
logic        cpu_data_we;
logic [31:0] cpu_data_addr;
logic [31:0] cpu_data_wdata;
logic [31:0] cpu_data_rdata;

//data sram
logic        data_sram_en;
logic        data_sram_we;
logic [31:0] data_sram_addr;
logic [31:0] data_sram_wdata;
logic [31:0] data_sram_rdata;

//conf
logic        conf_en;
logic        conf_we;
logic [31:0] conf_addr;
logic [31:0] conf_wdata;
logic [31:0] conf_rdata;
logic [15:0] conf_led;

//cpu
minicpu_top cpu(
    .clk              (cpu_clk       ),
    .resetn           (cpu_resetn    ),  //low active

    .inst_sram_we     (cpu_inst_we   ),
    .inst_sram_addr   (cpu_inst_addr ),
    .inst_sram_wdata  (cpu_inst_wdata),
    .inst_sram_rdata  (cpu_inst_rdata),
   
    .data_sram_we     (cpu_data_we   ),
    .data_sram_addr   (cpu_data_addr ),
    .data_sram_wdata  (cpu_data_wdata),
    .data_sram_rdata  (cpu_data_rdata)
);

assign cpu_data_rdata = (cpu_data_addr == 32'd1024)? {24'b0, ~switch_1[7:0]} :
                                                      32'b0;

//inst ram
inst_ram inst_ram
(
    .clk   (cpu_clk            ),   
    .we    (cpu_inst_we        ),   
    .a     (cpu_inst_addr[16:2]),   
    .d     (cpu_inst_wdata     ),   
    .spo   (cpu_inst_rdata     )   
);

//confreg
confreg u_confreg
(
    .clk          ( cpu_clk    ),  // i, 1   
    .resetn       ( cpu_resetn ),  // i, 1    
    .conf_we      ( conf_we    ),  // i, 4      
    .conf_wdata   ( conf_wdata ),  // i, 32         
    .led          ( conf_led   )   // o, 16   
);

assign conf_we    = cpu_data_we && cpu_data_addr == 32'd1028;
assign conf_wdata = cpu_data_wdata;

assign led = ~conf_led; 

endmodule

